module tb_regfile(output err);
  // your implementation here
endmodule: tb_regfile
