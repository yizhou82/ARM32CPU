module tb_datapath(output err);
  // your implementation here
endmodule: tb_datapath
