module tb_idecoder(output err);

endmodule: tb_idecoder