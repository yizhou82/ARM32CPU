module tb_ALU(output err);
  // your implementation here
endmodule: tb_ALU
