module tb_shifter(output err);
  // your implementation here
endmodule: tb_shifter
